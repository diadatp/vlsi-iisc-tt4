`default_nettype none

module note_lut (
    input clk,
    input rstn,
    input [3:0] note,
    input [3:0] octave,
    output reg [15:0] div
);

  reg [15:0] div_pre;

  // the lut is formed by assuming a clock frequency of 1MHz
  // div is the clock dividier required to geenrate the required frequency
  // divs = [int(1e6 / (16.35 * (2**(i / 12)))) for i in range(12)]
  // print("\n".join(divs)) <- not working TODO

  always @(posedge clk) begin
    case (note)
      4'h0: div_pre = 16'd61162;
      4'h1: div_pre = 16'd57729;
      4'h2: div_pre = 16'd54489;
      4'h3: div_pre = 16'd51430;
      4'h4: div_pre = 16'd48544;
      4'h5: div_pre = 16'd45819;
      4'h6: div_pre = 16'd43248;
      4'h7: div_pre = 16'd40820;
      4'h8: div_pre = 16'd38529;
      4'h9: div_pre = 16'd36367;
      4'hA: div_pre = 16'd34326;
      4'hB: div_pre = 16'd32399;
      default: div_pre = 16'd3822;
    endcase
  end

  always @(posedge clk) begin
    case (octave)
      4'd0: div = div_pre >> 0;
      4'd1: div = div_pre >> 1;
      4'd2: div = div_pre >> 2;
      4'd3: div = div_pre >> 3;
      4'd4: div = div_pre >> 4;
      4'd5: div = div_pre >> 5;
      4'd6: div = div_pre >> 6;
      4'd7: div = div_pre >> 7;
      4'd8: div = div_pre >> 8;
      default: div = div_pre;
    endcase
  end

endmodule
